// ECE:3350 SISC computer project
// finite state machine

`timescale 1ns/100ps


//TODO: Add the additional 6 internal signals to the parameter list
module ctrl (clk, rst_f, opcode, mm, stat, rf_we, alu_op, wb_sel, RB_SEL, BR_SEL, PC_RST, PC_WRITE, PC_SEL, IR_LOAD);

  /* TODO: Declare the additional internal signals listed above as inputs or outputs */
  
  input clk, rst_f;
  input [3:0] opcode, mm, stat;
  output reg rf_we,RB_SEL, BR_SEL, PC_RST, PC_WRITE, PC_SEL, IR_LOAD,wb_sel;
  output reg [1:0] alu_op;
  
  
  // state parameter declarations
  parameter start0 = 0, start1 = 1, fetch = 2, decode = 3, execute = 4, mem = 5, writeback = 6;
   
  // opcode paramenter declarations
  parameter NOOP = 0, LOD = 1, STR = 2, SWP = 3, BRA = 4, BRR = 5, BNE = 6, BNR = 7, ALU_OP = 8, HLT=15;

  // addressing modes
  parameter AM_IMM = 8;

  // state register and next state value
  reg [2:0]  present_state, next_state;

  // Initialize present state to 'start0'.
  initial
    present_state = start0;

  /* Clock procedure that progresses the fsm to the next state on the positive 
     edge of the clock, OR resets the state to 'start1' on the negative edge
     of rst_f. Notice that the computer is reset when rst_f is low, not high. */

  always @(posedge clk, negedge rst_f)
  begin
    if (rst_f == 1'b0)
      present_state <= start1;
    else
      present_state <= next_state;
  end
  
  /* Combinational procedure that determines the next state of the fsm. */

  always @(present_state, rst_f)
  begin
    case(present_state)
      start0:
        next_state = start1;
      start1:
	if (rst_f == 1'b0) 
          next_state = start1;
	else
          next_state = fetch;
      fetch:
        next_state = decode;
      decode:
        next_state = execute;
      execute:
        next_state = mem;
      mem:
        next_state = writeback;
      writeback:
        next_state = fetch;
      default:
        next_state = start1;
    endcase
  end
  



  always @(present_state, opcode, mm)
  begin

  /* TODO: Put your default assignments for the additional 6 internal signals here.  */
    rf_we  = 1'b0;
    wb_sel = 1'b0;
    alu_op = 2'b10;
    RB_SEL = 1'b0;
    BR_SEL = 1'b0;
    PC_RST = 1'b0; 
    PC_WRITE = 1'b0; 
    PC_SEL = 1'b0;
    IR_LOAD = 1'b0; 
  
    case(present_state)
     start1:
      begin
        /*TODO: Set PC_RST*/
	PC_RST = 1'b1;
	
      end

      fetch:
      begin
        /*TODO: Set IR_LOAD and PC_WRITE*/
	IR_LOAD = 1'b1;
	PC_WRITE = 1'b1;
      end

      decode:
      begin
        /*TODO: Set PC_SEL and set BR_SEL and PC_WRITE based on different instructions*/
	PC_WRITE = 1'b0;
	
	if (opcode == BRA)
		begin
		if((mm & stat) != 0)
			begin
			PC_SEL = 1'b1; 
			BR_SEL = 1'b1;
			PC_WRITE = 1'b1;
			end
		end
	if (opcode == BRR)
		begin
		if((mm & stat) != 0)
			begin
			PC_SEL = 1'b1;
			BR_SEL = 1'b0;
			PC_WRITE = 1'b1;
			end
		end
	if (opcode == BNR)
		begin
		if((mm & stat) == 0)
			begin
			PC_SEL = 1'b1;
			BR_SEL = 1'b0;
			PC_WRITE = 1'b1;
			end
		end
	if (opcode == BNE)
		begin
		if((mm & stat) == 0)
			begin
			PC_SEL = 1'b1;
			BR_SEL = 1'b1;
			PC_WRITE = 1'b1;
			end
		end
      end

      execute:
      begin
        if ((opcode == ALU_OP) && (mm == AM_IMM))
          alu_op = 2'b01;
        else
          alu_op = 2'b00;
      end

      mem:
      begin
        if ((opcode == ALU_OP) && (mm == AM_IMM))
          alu_op = 2'b11;
        else
          alu_op = 2'b10;
      end

      writeback:
      begin
        if (opcode == ALU_OP)
          rf_we = 1'b1;  
      end

      default:
      begin
      
      /* TODO: Put your default assignments for the additional 6 internal signals here.  */
        rf_we  = 1'b0;
        wb_sel = 1'b0;
        alu_op = 2'b10;
  	RB_SEL = 1'b0;
    	BR_SEL = 1'b0;
    	PC_RST = 1'b0;
    	PC_WRITE = 1'b0;
    	PC_SEL = 1'b0;
    	IR_LOAD = 1'b0;
      end
    endcase
  end

// Halt on HLT instruction  
  always @(opcode)
  begin
    if (opcode == HLT)
    begin 
      #5 $display ("Halt."); //Delay 5 ns so $monitor will print the halt instruction
      $stop;
    end
  end
    
  
endmodule
